`timescale 1ns/1ns
module test_cpu();
  reg clk, rst;
  always #100 clk = ~clk;
  CPU c(clk, rst);
  
  initial begin
   clk = 0 ;
   rst = 1 ;
   #500 ;
   rst =0 ;
   #4200 ;
   $stop ;
  end
endmodule

